// A clock that outputs 1 every n ticks.
mod clock(period) {
    let n = n + 1;
    output((n % period) == 0);
}

// A register that stores a single value.
mod cell(clk,write,val) {
    let stored = clk & write ? val : stored;
    output(stored);
}

// Converts a digit into signals to drive a 7 segment display.
// Compiled as a separate blueprint.
mod segments(x: $X) -> ($A,$B,$C,$D,$E,$F,$G) {

    let y = match(x) {
        0 => 0b0111111,
        1 => 6,
        2 => 91,
        3 => 79,
        4 => 102,
        5 => 109,
        6 => 125,
        7 => 0b0000111,
        8 => 0b1111111,
        9 => 111
    };

    output(y&1, y&2, y&4, y&8, y&16, y&32, y&64);
}

mod sqrt_step(S,x) {
    output((S/x + x)/2);
}

mod main(S) {
    let clk = clock(10);
    let val = cell(clk,1,next);
    let next = sqrt_step(S,val > 0 ? +val : 1);

    output(next);
}













/*
mod gpu_slice(C_Y,clk,data,y,write,clear) {
    let row_selected = C_Y == y;
    let $stored = 0;
    let new_val = stored ^ data;
    let $stored = cell(clk,write & row_selected,new_val);
    let collision = if(row_selected, new_val < stored, 0);
    output(stored); // new_val < stored
}

mod main(data,x,y,write,clear) {
    let clk = clock(30);

    let write_low = write & (x < 32);
    let data_low = data << x;

    let r0 = gpu_slice(0,    clk,data_low,y,write_low,clear);
    let r1 = gpu_slice(1,    clk,data_low,y,write_low,clear);
    let r2 = gpu_slice(2,    clk,data_low,y,write_low,clear);
    let r3 = gpu_slice(3,    clk,data_low,y,write_low,clear);
    output(r0,r1,r2,r3);
}

/*mod meme(x) {
    output(
        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +

        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +

        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +

        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +

        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +

        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +

        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +

        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +

        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +

        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x
    );
}*/
