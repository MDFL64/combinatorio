const MASK_ALU = 0xF;
    const ALU_ARG2  = 0x0;
    const ALU_OR    = 0x1;
    const ALU_AND   = 0x2;
    const ALU_XOR   = 0x3;
    const ALU_ADD   = 0x4;
    const ALU_SUB   = 0x5;
    const ALU_UP    = 0x6; // shift X up by 1
    const ALU_SUB2  = 0x7; // Y - X
    const ALU_EQ    = 0x8; // Not masked from 8XY* instruction
    const ALU_NEQ   = 0x9; // Not masked from 8XY* instruction
    const ALU_SPITE_ADDR = 0xA; // Not masked from 8XY* instruction
    const ALU_ARG1  = 0xB; // Not masked from 8XY* instruction
    const ALU_DOWN  = 0xE; // shift X down by 1

const MASK_PC = 0xF0;
    const PC_NEXT           = 0x00; // pc + 2
    const PC_GOTO           = 0x10; // res
    const PC_COND_SKIP      = 0x20; // res ? pc+4 : pc+2
    const PC_POP            = 0x30; // stack pop

const MASK_ARG1 = 0xF00;
    const ARG1_VX   = 0x000;
    const ARG1_RAND = 0x100;
    const ARG1_V0   = 0x200;

const MASK_ARG2 = 0xF000;
    const ARG2_VY           = 0x0000;
    const ARG2_IMM_8        = 0x1000;
    const ARG2_IMM_12       = 0x2000;
    const ARG2_KEY          = 0x3000;
    const ARG2_DELAY        = 0x4000;
    const ARG2_I            = 0x5000;

const MASK_WRITE = 0xF0000;
    const WRITE_VX      = 0x10000;
    const WRITE_I       = 0x20000;
    const WRITE_DELAY   = 0x30000;
    const WRITE_SOUND   = 0x40000;
    const WRITE_PUSH    = 0x50000; // write pc(+2?) to stack, sp++
    const WRITE_POP     = 0x60000; // sp--
    const WRITE_SCREEN  = 0x70000;
    const WRITE_CLS     = 0x80000;

const FLAG_STAY = 0x100000;

// ---- 00E0 = TODO clear screen
// 00EE = PC_POP | WRITE_POP
// 1NNN = PC_GOTO | ARG2_IMM_12
// 2NNN = PC_GOTO | ARG2_IMM_12 | WRITE_PUSH
// 3XNN = ALU_EQ | ARG2_IMM_8 | PC_COND_SKIP
// 4XNN = ALU_NEQ | ARG2_IMM_8 | PC_COND_SKIP
// 5XY0 = ALU_EQ | PC_COND_SKIP
// 6XNN = WRITE_VX | ARG2_IMM_8
// 7XNN = WRITE_VX | ALU_ADD | ARG2_IMM_8
// 8XYN = WRITE_VX | (instr & 0xF)
// 9XY0 = ALU_NEQ | PC_COND_SKIP
// ANNN = WRITE_I | ARG2_IMM_12
// BNNN = PC_GOTO | ALU_ADD | ARG1_V0 | ARG2_IMM_12
// CXNN = WRITE_VX | ALU_AND | ARG1_RAND | ARG2_IMM_8
// ---- DXYN = TODO draw sprite
// EX9E = ALU_EQ | PC_COND_SKIP | ARG2_KEY
// EXA1 = ALU_NEQ | PC_COND_SKIP | ARG2_KEY
// FX07 = WRITE_VX | ARG2_DELAY
// ---- FX0A = WRITE_VX | ARG2_KEY // TODO BLOCKS
// FX15 = WRITE_DELAY | ALU_ARG1
// FX18 = WRITE_SOUND | ALU_ARG1
// FX1E = WRITE_I | ALU_ADD | ARG2_I;
// FX29 = WRITE_I | ALU_SPRITE_ADDR
// ---- FX33 = TODO BCD
// ---- FX55 = TODO REG DUMP
// ---- FX65 = TODO REG LOAD


// Fibonacci
/*
mod rom(addr) {
    output(match(addr) {
        0 => 0x60, 1 => 0x00, // V0 = 0
        2 => 0x61, 3 => 0x01, // V1 = 1

        4 => 0x83, 5 => 0x00, // V3 = V0
        6 => 0x83, 7 => 0x14, // V3 = V3 + V1
        8 => 0x80, 9 => 0x10, // V0 = V1
        10 => 0x81, 11 => 0x30, // V1 = V3
        12 => 0x10, 13 => 0x04, // goto 004
    })
}*/

mod rom(addr) {
    output(match(addr) {
        0 => 0xA0, 1 => 20, // I = 20
        2 => 0x61, 3 => 0x00, // V1 = 0

        4 => 0x00, 5 => 0xE0, // cls

        6 => 0x60, 7 => 1, // V0 = 1
        8 => 0xD0, 9 => 0x18, // Draw @ (V0,V1)

        10 => 0x60, 11 => 8, // V0 = 10
        12 => 0xD0, 13 => 0x18, // Draw @ (V0,V1)

        14 => 0x60, 15 => 15, // V0 = 19
        16 => 0xD0, 17 => 0x18, // Draw @ (V0,V1)

        18 => 0x10, 19 => 0x04, // goto 04

        20 => 0x7e,     // sprite
        21 => 0x81,     // sprite
        22 => 0xa5,     // sprite
        23 => 0xa5,     // sprite
        24 => 0x81,     // sprite
        25 => 0xbd,     // sprite
        26 => 0x81,     // sprite
        27 => 0x7e,     // sprite
    });
}

mod decoder(instr,step) {
    let count = instr & 0xF;
    let cv = step < 1 ? FLAG_STAY : match(instr >> 12) {
        0 => match(instr) {
            0x00E0 => WRITE_CLS
        },
        1 => PC_GOTO | ARG2_IMM_12,
        6 => WRITE_VX | ARG2_IMM_8,
        7 => WRITE_VX | ALU_ADD | ARG2_IMM_8,
        8 => WRITE_VX | (instr & 0xF),
        0xA => WRITE_I | ALU_ARG2 | ARG2_IMM_12,
        0xD =>
            step==1 ? FLAG_STAY :
            step<count+1 ? WRITE_SCREEN | FLAG_STAY :
                WRITE_SCREEN
    };

    output(cv);
}

mod value_registers(x, y, write, write_val, clk) {
    let write_val_byte = write_val & 0xFF;
    let V0 = cell(clk,(x==0) & write,write_val_byte);
    let V1 = cell(clk,(x==1) & write,write_val_byte);
    let V2 = cell(clk,(x==2) & write,write_val_byte);
    let V3 = cell(clk,(x==3) & write,write_val_byte);
    let V4 = cell(clk,(x==4) & write,write_val_byte);
    let V5 = cell(clk,(x==5) & write,write_val_byte);
    let V6 = cell(clk,(x==6) & write,write_val_byte);
    let V7 = cell(clk,(x==7) & write,write_val_byte);
    let V8 = cell(clk,(x==8) & write,write_val_byte);
    let V9 = cell(clk,(x==9) & write,write_val_byte);
    let VA = cell(clk,(x==10) & write,write_val_byte);
    let VB = cell(clk,(x==11) & write,write_val_byte);
    let VC = cell(clk,(x==12) & write,write_val_byte);
    let VD = cell(clk,(x==13) & write,write_val_byte);
    let VE = cell(clk,(x==14) & write,write_val_byte);
    let VF = cell(clk,(x==15) & write,write_val_byte); // TODO specialized write to carry flag

    let res_x = match(x) {
        0 => V0,
        1 => V1,
        2 => V2,
        3 => V3,
        4 => V4,
        5 => V5,
        6 => V6,
        7 => V7,
        8 => V8,
        9 => V9,
        10 => VA,
        11 => VB,
        12 => VC,
        13 => VD,
        14 => VE,
        15 => VF
    };

    let res_y = match(y) {
        0 => V0,
        1 => V1,
        2 => V2,
        3 => V3,
        4 => V4,
        5 => V5,
        6 => V6,
        7 => V7,
        8 => V8,
        9 => V9,
        10 => VA,
        11 => VB,
        12 => VC,
        13 => VD,
        14 => VE,
        15 => VF
    };

    output(+res_x,+res_y,V0);
}

mod main(reset) -> ($DOT,$X,$Y,$D,$W,$C) {
    let clk = clock(30);

    let next_step = advance_instr ? 0 : step+1;
    let step = cell(clk,1,next_step);
    let pc = cell(clk,advance_instr,next_pc);
    let I = cell(clk,write_to_i,res & 0xFFF);

    let mem_read_addr = (step <= 1) ? (pc + step) : (I + step - 2);
    let mem_read_val = rom(mem_read_addr);

    // Current instruction
    let ir = cell(clk,1,instr);
    let instr = match(step) {
        0 => mem_read_val<<8,
        1 => ir | mem_read_val,
        >1 => ir
    };


    // The decoder gives us back a control vector
    let cv = decoder(instr,step);

    let advance_instr = !(cv & FLAG_STAY) | reset;
    
    let pc_inc = pc+2;
    let next_pc = reset ? 0 : match(cv & MASK_PC) {
        PC_NEXT => pc_inc,
        PC_GOTO => +res,
        PC_COND_SKIP => (res != 0) ? pc+4 : pc_inc,
        PC_POP => 0 // TODO
    };

    let write_select = cv & MASK_WRITE;
    let write_to_vx = write_select == WRITE_VX;
    let write_to_i = write_select == WRITE_I;
    let write_to_screen = write_select == WRITE_SCREEN;
    let clear_screen = write_select == WRITE_CLS;

    let x = (instr >> 8) & 0xF;
    let y = (instr >> 4) & 0xF;
    let (vx,vy,v0) = value_registers(x,y,write_to_vx,res,clk);

    let arg1 = vx;

    let arg2 = match(cv & MASK_ARG2) {
        ARG2_VY => vy,
        ARG2_IMM_8 => instr & 0xFF,
        ARG2_IMM_12 => instr & 0xFFF
    };

    let res = match(cv & MASK_ALU) {
        ALU_ARG2 => arg2,
        ALU_ADD => arg1 + arg2,
    };

    output(clk,vx,vy + (step-2),mem_read_val,write_to_screen,clear_screen)
}
