//use "std/math";

// Iteratively computes the square root of a positive integer.
// Takes time to run and likely can be optimized.
mod sqrt(S) {
    let clk = clock(3); // seems stable
    let stored = cell(clk,1,next);
    let x = max(stored,1); // get rid of negative values
    let next = (S/x + x)/2;
    output(next);
}

mod main(y) {
    output(123)
}

mod main(x) {
    output(clamp(1,abs(x),10));
}

// Converts a digit into signals to drive a 7 segment display.
// Compiled as a separate blueprint.
/*mod segments(x: $X) -> ($A,$B,$C,$D,$E,$F,$G) {

    let y = match(x) {
        0 => 0b0111111,
        1 => 0b0000110,
        2 => 0b1011011,
        3 => 0b1001111,
        4 => 0b1100110,
        5 => 0b1101101,
        6 => 0b1111101,
        7 => 0b0000111,
        8 => 0b1111111,
        9 => 0b1101111
    };

    output(y&1, y&2, y&4, y&8, y&16, y&32, y&64);
}*/









/*
mod gpu_slice(C_Y,clk,data,y,write,clear) {
    let row_selected = C_Y == y;
    let $stored = 0;
    let new_val = stored ^ data;
    let $stored = cell(clk,write & row_selected,new_val);
    let collision = if(row_selected, new_val < stored, 0);
    output(stored); // new_val < stored
}

mod main(data,x,y,write,clear) {
    let clk = clock(30);

    let write_low = write & (x < 32);
    let data_low = data << x;

    let r0 = gpu_slice(0,    clk,data_low,y,write_low,clear);
    let r1 = gpu_slice(1,    clk,data_low,y,write_low,clear);
    let r2 = gpu_slice(2,    clk,data_low,y,write_low,clear);
    let r3 = gpu_slice(3,    clk,data_low,y,write_low,clear);
    output(r0,r1,r2,r3);
}

/*mod meme(x) {
    output(
        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +

        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +

        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +

        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +

        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +

        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +

        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +

        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +

        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +

        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x +
        x+x+x+x+x+x+x+x+x+x
    );
}*/
